/* Module Name	: ECRC                      */
/* Written By	: Mohamed Khaled Alahmady   */
/* Date			: 29-04-2024		        */
/* Version		: V_1			            */
/* Updates		: -			                */
/* Dependencies	: -				            */
/* Used			: -			                */
module ECRC #(
)(
	input bit clk,
    input bit arst,
    // Interface with Fragmentation
    Fragmentation_Interface.ECRC_FRAGMENTATION   _if
);

/* Packages */
import Fragmentation_Package::*;

/* Parameters */

/* Useful Functions */

/* Internal Signals */
reg [ECRC_POLY_WIDTH - 1 : 0] temp_seed;

/* Assign Statements */

/* Always Blocks */
always_ff @(posedge clk or negedge arst) begin
	if (!arst) begin
		_if.ecrc_Result_reg		<= '0;
	end
	else begin
		if(_if.ecrc_EN)
			_if.ecrc_Result_reg	<= _if.ecrc_Result_comb;		
	end
end

always @(*) begin
    if (_if.ecrc_EN) begin
		temp_seed = (_if.ecrc_Seed_Load) ? _if.ecrc_Seed : _if.ecrc_Result_reg;
        // Data Length 32 bits	(1DW)
		if (_if.ecrc_Length == 'd1) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[  0] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 17] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 18] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[  0] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 29]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 28]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 27]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 26]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[  0] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 10] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 11] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 12] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 28]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 27]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26]);
		end		
        // Data Length 64 bits	(2DW)
		else if (_if.ecrc_Length == 'd2) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 12] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 13] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[  0] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 61]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 60]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 59]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 58]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[  0] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[  1] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 61]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[  2] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 60]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 59]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 58]);
		end	
        // Data Length 96 bits	(3DW)
		else if (_if.ecrc_Length == 'd3) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 23] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 95]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[  0] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 93]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 92]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 91]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 90]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 95]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 94]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[  0] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 93]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 92]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 91]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 90]);
		end	
		// Data Length 128 bits	(4DW)
		else if (_if.ecrc_Length == 'd4) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[127]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[125]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[124]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[123]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[122]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[127]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 40] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 90] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[125]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 39] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 54] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 89] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[127]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 38] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 53] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 88] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[126]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[  8] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 21] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 37] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 52] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 59] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 87] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[125]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  7] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 20] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 36] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 51] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 58] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 72] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 77] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 86] ^ _if.ecrc_Message[ 93] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[124]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  4] ^ _if.ecrc_Message[  6] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 13] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 16] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 19] ^ _if.ecrc_Message[ 23] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 26] ^ _if.ecrc_Message[ 28] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 35] ^ _if.ecrc_Message[ 42] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 48] ^ _if.ecrc_Message[ 50] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 57] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 64] ^ _if.ecrc_Message[ 66] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 69] ^ _if.ecrc_Message[ 71] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 76] ^ _if.ecrc_Message[ 79] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 82] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 85] ^ _if.ecrc_Message[ 92] ^ _if.ecrc_Message[ 95] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[123]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ _if.ecrc_Message[  0] ^ _if.ecrc_Message[  1] ^ _if.ecrc_Message[  2] ^ _if.ecrc_Message[  3] ^ _if.ecrc_Message[  5] ^ _if.ecrc_Message[  9] ^ _if.ecrc_Message[ 10] ^ _if.ecrc_Message[ 11] ^ _if.ecrc_Message[ 12] ^ _if.ecrc_Message[ 14] ^ _if.ecrc_Message[ 15] ^ _if.ecrc_Message[ 17] ^ _if.ecrc_Message[ 18] ^ _if.ecrc_Message[ 22] ^ _if.ecrc_Message[ 24] ^ _if.ecrc_Message[ 25] ^ _if.ecrc_Message[ 27] ^ _if.ecrc_Message[ 29] ^ _if.ecrc_Message[ 30] ^ _if.ecrc_Message[ 31] ^ _if.ecrc_Message[ 32] ^ _if.ecrc_Message[ 33] ^ _if.ecrc_Message[ 34] ^ _if.ecrc_Message[ 41] ^ _if.ecrc_Message[ 43] ^ _if.ecrc_Message[ 44] ^ _if.ecrc_Message[ 45] ^ _if.ecrc_Message[ 46] ^ _if.ecrc_Message[ 47] ^ _if.ecrc_Message[ 49] ^ _if.ecrc_Message[ 55] ^ _if.ecrc_Message[ 56] ^ _if.ecrc_Message[ 60] ^ _if.ecrc_Message[ 61] ^ _if.ecrc_Message[ 62] ^ _if.ecrc_Message[ 63] ^ _if.ecrc_Message[ 65] ^ _if.ecrc_Message[ 67] ^ _if.ecrc_Message[ 68] ^ _if.ecrc_Message[ 70] ^ _if.ecrc_Message[ 73] ^ _if.ecrc_Message[ 74] ^ _if.ecrc_Message[ 75] ^ _if.ecrc_Message[ 78] ^ _if.ecrc_Message[ 80] ^ _if.ecrc_Message[ 81] ^ _if.ecrc_Message[ 83] ^ _if.ecrc_Message[ 84] ^ _if.ecrc_Message[ 91] ^ _if.ecrc_Message[ 94] ^ _if.ecrc_Message[ 96] ^ _if.ecrc_Message[ 97] ^ _if.ecrc_Message[ 98] ^ _if.ecrc_Message[ 99] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[122]);
		end
		// Data Length 160 bits (5DW)
		else if (_if.ecrc_Length == 'd5) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[2] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[0] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[28] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[31] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[3] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2]);
		end	
        // Data Length 192 bits	(6DW)
		else if (_if.ecrc_Length == 'd6) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[6] 	^ temp_seed[7]  ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[6] 	^ temp_seed[8]  ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] 	^ temp_seed[6]  ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] 	^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[3] ^ temp_seed[7] ^ temp_seed[8] 	^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[4] 	^ temp_seed[6]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] 	^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] 	^ temp_seed[7]  ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] 	^ temp_seed[3]  ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] 	^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] 	^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[5] 	^ temp_seed[7]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[30] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[2] ^ temp_seed[5] ^ temp_seed[7] 	^ temp_seed[8]  ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[3] ^ temp_seed[6] ^ temp_seed[8] 	^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[7] 	^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5] 	^ temp_seed[8]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[0] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[1] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[2] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[31] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4]  ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2]  ^ temp_seed[5]  ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[3] ^ temp_seed[7] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2]  ^ temp_seed[4]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[31] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2]  ^ temp_seed[3]  ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3]  ^ temp_seed[4]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3]  ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[31] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[6]  ^ temp_seed[7]  ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[7]  ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5]  ^ temp_seed[6]  ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
		end	
        // Data Length 224 bits	(7DW)
		else if (_if.ecrc_Length == 'd7) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^_if.ecrc_Message[223] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[3] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9]  ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^_if.ecrc_Message[223] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[1] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5] ^ temp_seed[7]  ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[3] ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[8]  ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[2] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9]  ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[7]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[8]  ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[9]  ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[30] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[31] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[6]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[30] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[31] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[0]);
		end	
        // Data Length 256 bits	(8DW)
		else if (_if.ecrc_Length == 'd8) begin
			_if.ecrc_Result_comb[ 7] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[19] ^ temp_seed[24] ^ temp_seed[28] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 6] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 5] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 4] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 3] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[30] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 2] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4]);
			_if.ecrc_Result_comb[ 1] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[ 0] = ~(temp_seed[0] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[15] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[14] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[13] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5]);
			_if.ecrc_Result_comb[12] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[11] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[10] = ~(temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[ 9] = ~(temp_seed[0] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[ 8] = ~(temp_seed[1] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[30] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1]);
			
			_if.ecrc_Result_comb[23] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5]);
			_if.ecrc_Result_comb[22] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4]);
			_if.ecrc_Result_comb[21] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[20] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[19] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[18] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[17] = ~(temp_seed[1] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[83] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2]);
			_if.ecrc_Result_comb[16] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[30] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[82] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[1] ^ _if.ecrc_Message[0]);
			
			_if.ecrc_Result_comb[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[31] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[239] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[81] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[39] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[30] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[238] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[218] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[168] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[80] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[38] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[3]);
			_if.ecrc_Result_comb[29] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[13] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[255] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[237] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[217] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[182] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[167] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[118] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[79] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[37] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[18] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[28] = ~(temp_seed[1] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[254] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[236] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[216] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[181] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[166] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[117] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[111] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[78] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[36] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[17] ^ _if.ecrc_Message[12] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[27] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[253] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[243] ^ _if.ecrc_Message[235] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[215] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[187] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[180] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[165] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[149] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[136] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[127] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[116] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[110] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[104] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[93] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[77] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[52] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[35] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[25] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[16] ^ _if.ecrc_Message[11] ^ _if.ecrc_Message[7] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[26] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[30] ^ _if.ecrc_Message[252] ^ _if.ecrc_Message[249] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[242] ^ _if.ecrc_Message[234] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[221] ^ _if.ecrc_Message[214] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[205] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[200] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[186] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[179] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[164] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[148] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[135] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[126] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[115] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[109] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[103] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[97] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[92] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[76] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[72] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[61] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[51] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[34] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[24] ^ _if.ecrc_Message[21] ^ _if.ecrc_Message[15] ^ _if.ecrc_Message[10] ^ _if.ecrc_Message[6] ^ _if.ecrc_Message[3] ^ _if.ecrc_Message[1]);
			_if.ecrc_Result_comb[25] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[17] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[31] ^ _if.ecrc_Message[251] ^ _if.ecrc_Message[248] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[245] ^ _if.ecrc_Message[241] ^ _if.ecrc_Message[233] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[229] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[223] ^ _if.ecrc_Message[220] ^ _if.ecrc_Message[213] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[210] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[207] ^ _if.ecrc_Message[204] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[199] ^ _if.ecrc_Message[197] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[194] ^ _if.ecrc_Message[192] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[185] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[178] ^ _if.ecrc_Message[176] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[170] ^ _if.ecrc_Message[163] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[156] ^ _if.ecrc_Message[154] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[151] ^ _if.ecrc_Message[147] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[144] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[141] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[134] ^ _if.ecrc_Message[132] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[125] ^ _if.ecrc_Message[123] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[114] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[108] ^ _if.ecrc_Message[106] ^ _if.ecrc_Message[102] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[99] ^ _if.ecrc_Message[96] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[91] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[88] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[75] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[71] ^ _if.ecrc_Message[69] ^ _if.ecrc_Message[67] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[60] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[56] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[50] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[45] ^ _if.ecrc_Message[43] ^ _if.ecrc_Message[41] ^ _if.ecrc_Message[33] ^ _if.ecrc_Message[31] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[27] ^ _if.ecrc_Message[23] ^ _if.ecrc_Message[20] ^ _if.ecrc_Message[14] ^ _if.ecrc_Message[9] ^ _if.ecrc_Message[5] ^ _if.ecrc_Message[2] ^ _if.ecrc_Message[0]);
			_if.ecrc_Result_comb[24] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[18] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[30] ^ _if.ecrc_Message[250] ^ _if.ecrc_Message[247] ^ _if.ecrc_Message[246] ^ _if.ecrc_Message[244] ^ _if.ecrc_Message[240] ^ _if.ecrc_Message[232] ^ _if.ecrc_Message[231] ^ _if.ecrc_Message[230] ^ _if.ecrc_Message[228] ^ _if.ecrc_Message[227] ^ _if.ecrc_Message[226] ^ _if.ecrc_Message[225] ^ _if.ecrc_Message[224] ^ _if.ecrc_Message[222] ^ _if.ecrc_Message[219] ^ _if.ecrc_Message[212] ^ _if.ecrc_Message[211] ^ _if.ecrc_Message[209] ^ _if.ecrc_Message[208] ^ _if.ecrc_Message[206] ^ _if.ecrc_Message[203] ^ _if.ecrc_Message[202] ^ _if.ecrc_Message[201] ^ _if.ecrc_Message[198] ^ _if.ecrc_Message[196] ^ _if.ecrc_Message[195] ^ _if.ecrc_Message[193] ^ _if.ecrc_Message[191] ^ _if.ecrc_Message[190] ^ _if.ecrc_Message[189] ^ _if.ecrc_Message[188] ^ _if.ecrc_Message[184] ^ _if.ecrc_Message[183] ^ _if.ecrc_Message[177] ^ _if.ecrc_Message[175] ^ _if.ecrc_Message[174] ^ _if.ecrc_Message[173] ^ _if.ecrc_Message[172] ^ _if.ecrc_Message[171] ^ _if.ecrc_Message[169] ^ _if.ecrc_Message[162] ^ _if.ecrc_Message[161] ^ _if.ecrc_Message[160] ^ _if.ecrc_Message[159] ^ _if.ecrc_Message[158] ^ _if.ecrc_Message[157] ^ _if.ecrc_Message[155] ^ _if.ecrc_Message[153] ^ _if.ecrc_Message[152] ^ _if.ecrc_Message[150] ^ _if.ecrc_Message[146] ^ _if.ecrc_Message[145] ^ _if.ecrc_Message[143] ^ _if.ecrc_Message[142] ^ _if.ecrc_Message[140] ^ _if.ecrc_Message[139] ^ _if.ecrc_Message[138] ^ _if.ecrc_Message[137] ^ _if.ecrc_Message[133] ^ _if.ecrc_Message[131] ^ _if.ecrc_Message[130] ^ _if.ecrc_Message[129] ^ _if.ecrc_Message[128] ^ _if.ecrc_Message[124] ^ _if.ecrc_Message[122] ^ _if.ecrc_Message[121] ^ _if.ecrc_Message[120] ^ _if.ecrc_Message[119] ^ _if.ecrc_Message[113] ^ _if.ecrc_Message[112] ^ _if.ecrc_Message[107] ^ _if.ecrc_Message[105] ^ _if.ecrc_Message[101] ^ _if.ecrc_Message[100] ^ _if.ecrc_Message[98] ^ _if.ecrc_Message[95] ^ _if.ecrc_Message[94] ^ _if.ecrc_Message[90] ^ _if.ecrc_Message[89] ^ _if.ecrc_Message[87] ^ _if.ecrc_Message[86] ^ _if.ecrc_Message[85] ^ _if.ecrc_Message[84] ^ _if.ecrc_Message[74] ^ _if.ecrc_Message[73] ^ _if.ecrc_Message[70] ^ _if.ecrc_Message[68] ^ _if.ecrc_Message[66] ^ _if.ecrc_Message[65] ^ _if.ecrc_Message[64] ^ _if.ecrc_Message[63] ^ _if.ecrc_Message[62] ^ _if.ecrc_Message[59] ^ _if.ecrc_Message[58] ^ _if.ecrc_Message[57] ^ _if.ecrc_Message[55] ^ _if.ecrc_Message[54] ^ _if.ecrc_Message[53] ^ _if.ecrc_Message[49] ^ _if.ecrc_Message[48] ^ _if.ecrc_Message[47] ^ _if.ecrc_Message[46] ^ _if.ecrc_Message[44] ^ _if.ecrc_Message[42] ^ _if.ecrc_Message[40] ^ _if.ecrc_Message[32] ^ _if.ecrc_Message[30] ^ _if.ecrc_Message[29] ^ _if.ecrc_Message[28] ^ _if.ecrc_Message[26] ^ _if.ecrc_Message[22] ^ _if.ecrc_Message[19] ^ _if.ecrc_Message[13] ^ _if.ecrc_Message[8] ^ _if.ecrc_Message[4] ^ _if.ecrc_Message[1]);
		end	
        else begin
            _if.ecrc_Result_comb   = {ECRC_POLY_WIDTH{1'b0}};
        end
    end
    else begin
        _if.ecrc_Result_comb   = {ECRC_POLY_WIDTH{1'b0}};
    end
end

/* Instantiations */

endmodule: ECRC
/*********** END_OF_FILE ***********/