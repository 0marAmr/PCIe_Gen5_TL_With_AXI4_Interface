/* Module Name	: CRC32_Parallel				*/
/* Written By	: Ahmady                     	*/
/* Date			: 26-02-2024					*/
/* Version		: V_1							*/
/* Updates		: -								*/
/* Dependencies	: -								*/
/* Used			: - 							*/
/* Synthesizable: YES                           */
`timescale 1ns/1ps
module CRC32_Parallel #(
    parameter   DATA_WIDTH 		= 256,      // Data Bus Width (8DW from TL to DLL)
				LENGTH_WIDTH 	= 4,        // Length of Valid Data in DW
                POLY_WIDTH 		= 32        // Polynomial Order (for PCIe 32-bits 0x04C11DB7) 
)(
	input 	wire [DATA_WIDTH - 1 : 0]     	CRC_i_Message,
	input   wire [LENGTH_WIDTH - 1 : 0]   	CRC_i_Length,
	input 	wire                        	CRC_i_EN,	
    input   wire [POLY_WIDTH - 1 : 0]		CRC_i_Seed,             
    input   wire 							CRC_i_Seed_Load,    
	// Number of Cycles [8] bits
	output 	reg  [POLY_WIDTH - 1 : 0]   	CRC_o_CRC
);

/* Parameters (must be in upper case) */

/* Internal Signals */
reg [POLY_WIDTH - 1 : 0] temp_seed;

/* Assign Statements */

/* Always Blocks */
always @(*) begin
    if (CRC_i_EN) begin
		temp_seed = (CRC_i_Seed_Load) ? CRC_i_Seed : CRC_o_CRC;
        // Data Length 32 bits	(1DW)
		if (CRC_i_Length == 'd1) begin
			CRC_o_CRC[ 7] = ~(temp_seed[  0] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[ 6] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[ 5] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[ 4] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[ 3] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[ 2] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[ 1] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  6] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[ 0] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31]);
			
			CRC_o_CRC[15] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 17] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[14] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 18] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[13] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[12] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[11] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[10] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  6] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[ 9] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  5] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29]);
			CRC_o_CRC[ 8] = ~(temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28]);
			
			CRC_o_CRC[23] = ~(temp_seed[  0] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[22] = ~(temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[21] = ~(temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 29]);
			CRC_o_CRC[20] = ~(temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 28]);
			CRC_o_CRC[19] = ~(temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 27]);
			CRC_o_CRC[18] = ~(temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 26]);
			CRC_o_CRC[17] = ~(temp_seed[  0] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[16] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31]);
			
			CRC_o_CRC[31] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[30] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29]);
			CRC_o_CRC[29] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 10] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31]);
			CRC_o_CRC[28] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 11] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30]);
			CRC_o_CRC[27] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 12] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29]);
			CRC_o_CRC[26] = ~(temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 28]);
			CRC_o_CRC[25] = ~(temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 27]);
			CRC_o_CRC[24] = ~(temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26]);
		end		
        // Data Length 64 bits	(2DW)
		else if (CRC_i_Length == 'd2) begin
			CRC_o_CRC[ 7] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[ 6] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[ 5] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 12] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[ 4] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 13] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[ 3] = ~(temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[ 2] = ~(temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[ 1] = ~(temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[ 0] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63]);
			
			CRC_o_CRC[15] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[14] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[13] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[12] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[11] = ~(temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[10] = ~(temp_seed[  0] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[ 9] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61]);
			CRC_o_CRC[ 8] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60]);
			
			CRC_o_CRC[23] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[22] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[21] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 61]);
			CRC_o_CRC[20] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 60]);
			CRC_o_CRC[19] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 59]);
			CRC_o_CRC[18] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 58]);
			CRC_o_CRC[17] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[16] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63]);
			
			CRC_o_CRC[31] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[30] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61]);
			CRC_o_CRC[29] = ~(temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63]);
			CRC_o_CRC[28] = ~(temp_seed[  0] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62]);
			CRC_o_CRC[27] = ~(temp_seed[  1] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 61]);
			CRC_o_CRC[26] = ~(temp_seed[  2] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 60]);
			CRC_o_CRC[25] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 59]);
			CRC_o_CRC[24] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 58]);
		end	
        // Data Length 96 bits	(3DW)
		else if (CRC_i_Length == 'd3) begin
			CRC_o_CRC[ 7] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[ 6] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[ 5] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[ 4] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[ 3] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[ 2] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[ 1] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[ 0] = ~(temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 23] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 95]);
			
			CRC_o_CRC[15] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[14] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[13] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[12] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[11] = ~(temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[10] = ~(temp_seed[  0] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[ 9] = ~(temp_seed[  1] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93]);
			CRC_o_CRC[ 8] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92]);
			
			CRC_o_CRC[23] = ~(temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[22] = ~(temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[21] = ~(temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 93]);
			CRC_o_CRC[20] = ~(temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 92]);
			CRC_o_CRC[19] = ~(temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 91]);
			CRC_o_CRC[18] = ~(temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 90]);
			CRC_o_CRC[17] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 15] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[16] = ~(temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95]);
			
			CRC_o_CRC[31] = ~(temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[30] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93]);
			CRC_o_CRC[29] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 95]);
			CRC_o_CRC[28] = ~(temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 94]);
			CRC_o_CRC[27] = ~(temp_seed[  0] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 93]);
			CRC_o_CRC[26] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 92]);
			CRC_o_CRC[25] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 91]);
			CRC_o_CRC[24] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 90]);
		end	
		// Data Length 128 bits	(4DW)
		else if (CRC_i_Length == 'd4) begin
			CRC_o_CRC[ 7] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[111] ^ CRC_i_Message[115] ^ CRC_i_Message[117] ^ CRC_i_Message[118] ^ CRC_i_Message[121] ^ CRC_i_Message[127]);
			CRC_o_CRC[ 6] = ~(temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[103] ^ CRC_i_Message[110] ^ CRC_i_Message[111] ^ CRC_i_Message[114] ^ CRC_i_Message[115] ^ CRC_i_Message[116] ^ CRC_i_Message[118] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			CRC_o_CRC[ 5] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 97] ^ CRC_i_Message[101] ^ CRC_i_Message[103] ^ CRC_i_Message[109] ^ CRC_i_Message[110] ^ CRC_i_Message[111] ^ CRC_i_Message[113] ^ CRC_i_Message[114] ^ CRC_i_Message[118] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[125] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			CRC_o_CRC[ 4] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[100] ^ CRC_i_Message[102] ^ CRC_i_Message[108] ^ CRC_i_Message[109] ^ CRC_i_Message[110] ^ CRC_i_Message[112] ^ CRC_i_Message[113] ^ CRC_i_Message[117] ^ CRC_i_Message[118] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[124] ^ CRC_i_Message[125] ^ CRC_i_Message[126]);
			CRC_o_CRC[ 3] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 98] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[107] ^ CRC_i_Message[108] ^ CRC_i_Message[109] ^ CRC_i_Message[112] ^ CRC_i_Message[115] ^ CRC_i_Message[116] ^ CRC_i_Message[119] ^ CRC_i_Message[121] ^ CRC_i_Message[123] ^ CRC_i_Message[124] ^ CRC_i_Message[125] ^ CRC_i_Message[127]);
			CRC_o_CRC[ 2] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[103] ^ CRC_i_Message[106] ^ CRC_i_Message[107] ^ CRC_i_Message[108] ^ CRC_i_Message[114] ^ CRC_i_Message[117] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[124] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			CRC_o_CRC[ 1] = ~(temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 98] ^ CRC_i_Message[102] ^ CRC_i_Message[105] ^ CRC_i_Message[106] ^ CRC_i_Message[107] ^ CRC_i_Message[113] ^ CRC_i_Message[116] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[125] ^ CRC_i_Message[126]);
			CRC_o_CRC[ 0] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[105] ^ CRC_i_Message[106] ^ CRC_i_Message[111] ^ CRC_i_Message[112] ^ CRC_i_Message[117] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[122] ^ CRC_i_Message[124] ^ CRC_i_Message[125] ^ CRC_i_Message[127]);
			
			CRC_o_CRC[15] = ~(temp_seed[  1] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 99] ^ CRC_i_Message[104] ^ CRC_i_Message[105] ^ CRC_i_Message[110] ^ CRC_i_Message[115] ^ CRC_i_Message[116] ^ CRC_i_Message[117] ^ CRC_i_Message[119] ^ CRC_i_Message[123] ^ CRC_i_Message[124] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			CRC_o_CRC[14] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 98] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[109] ^ CRC_i_Message[114] ^ CRC_i_Message[115] ^ CRC_i_Message[116] ^ CRC_i_Message[118] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[125] ^ CRC_i_Message[126]);
			CRC_o_CRC[13] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[101] ^ CRC_i_Message[108] ^ CRC_i_Message[111] ^ CRC_i_Message[113] ^ CRC_i_Message[114] ^ CRC_i_Message[118] ^ CRC_i_Message[122] ^ CRC_i_Message[124] ^ CRC_i_Message[125] ^ CRC_i_Message[127]);
			CRC_o_CRC[12] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[107] ^ CRC_i_Message[110] ^ CRC_i_Message[111] ^ CRC_i_Message[112] ^ CRC_i_Message[113] ^ CRC_i_Message[115] ^ CRC_i_Message[118] ^ CRC_i_Message[123] ^ CRC_i_Message[124] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			CRC_o_CRC[11] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 97] ^ CRC_i_Message[100] ^ CRC_i_Message[103] ^ CRC_i_Message[106] ^ CRC_i_Message[109] ^ CRC_i_Message[110] ^ CRC_i_Message[112] ^ CRC_i_Message[114] ^ CRC_i_Message[115] ^ CRC_i_Message[118] ^ CRC_i_Message[121] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[125] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			CRC_o_CRC[10] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[ 10] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 99] ^ CRC_i_Message[102] ^ CRC_i_Message[105] ^ CRC_i_Message[108] ^ CRC_i_Message[109] ^ CRC_i_Message[111] ^ CRC_i_Message[113] ^ CRC_i_Message[114] ^ CRC_i_Message[117] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[122] ^ CRC_i_Message[124] ^ CRC_i_Message[125] ^ CRC_i_Message[126]);
			CRC_o_CRC[ 9] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 11] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 98] ^ CRC_i_Message[101] ^ CRC_i_Message[104] ^ CRC_i_Message[107] ^ CRC_i_Message[108] ^ CRC_i_Message[110] ^ CRC_i_Message[112] ^ CRC_i_Message[113] ^ CRC_i_Message[116] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[123] ^ CRC_i_Message[124] ^ CRC_i_Message[125]);
			CRC_o_CRC[ 8] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 97] ^ CRC_i_Message[100] ^ CRC_i_Message[103] ^ CRC_i_Message[106] ^ CRC_i_Message[107] ^ CRC_i_Message[109] ^ CRC_i_Message[111] ^ CRC_i_Message[112] ^ CRC_i_Message[115] ^ CRC_i_Message[118] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[124]);
			
			CRC_o_CRC[23] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 98] ^ CRC_i_Message[101] ^ CRC_i_Message[103] ^ CRC_i_Message[105] ^ CRC_i_Message[106] ^ CRC_i_Message[108] ^ CRC_i_Message[110] ^ CRC_i_Message[114] ^ CRC_i_Message[115] ^ CRC_i_Message[119] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[127]);
			CRC_o_CRC[22] = ~(temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 97] ^ CRC_i_Message[100] ^ CRC_i_Message[102] ^ CRC_i_Message[104] ^ CRC_i_Message[105] ^ CRC_i_Message[107] ^ CRC_i_Message[109] ^ CRC_i_Message[113] ^ CRC_i_Message[114] ^ CRC_i_Message[118] ^ CRC_i_Message[121] ^ CRC_i_Message[122] ^ CRC_i_Message[126]);
			CRC_o_CRC[21] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 99] ^ CRC_i_Message[101] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[106] ^ CRC_i_Message[108] ^ CRC_i_Message[112] ^ CRC_i_Message[113] ^ CRC_i_Message[117] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[125]);
			CRC_o_CRC[20] = ~(temp_seed[  1] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 98] ^ CRC_i_Message[100] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[105] ^ CRC_i_Message[107] ^ CRC_i_Message[111] ^ CRC_i_Message[112] ^ CRC_i_Message[116] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[124]);
			CRC_o_CRC[19] = ~(temp_seed[  2] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 99] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[104] ^ CRC_i_Message[106] ^ CRC_i_Message[110] ^ CRC_i_Message[111] ^ CRC_i_Message[115] ^ CRC_i_Message[118] ^ CRC_i_Message[119] ^ CRC_i_Message[123]);
			CRC_o_CRC[18] = ~(temp_seed[  0] ^ temp_seed[  3] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 98] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[103] ^ CRC_i_Message[105] ^ CRC_i_Message[109] ^ CRC_i_Message[110] ^ CRC_i_Message[114] ^ CRC_i_Message[117] ^ CRC_i_Message[118] ^ CRC_i_Message[122]);
			CRC_o_CRC[17] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 98] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[108] ^ CRC_i_Message[109] ^ CRC_i_Message[111] ^ CRC_i_Message[113] ^ CRC_i_Message[115] ^ CRC_i_Message[116] ^ CRC_i_Message[118] ^ CRC_i_Message[127]);
			CRC_o_CRC[16] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 98] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[107] ^ CRC_i_Message[108] ^ CRC_i_Message[110] ^ CRC_i_Message[111] ^ CRC_i_Message[112] ^ CRC_i_Message[114] ^ CRC_i_Message[118] ^ CRC_i_Message[121] ^ CRC_i_Message[126] ^ CRC_i_Message[127]);
			
			CRC_o_CRC[31] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 20] ^ temp_seed[ 22] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 29] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  2] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[106] ^ CRC_i_Message[107] ^ CRC_i_Message[109] ^ CRC_i_Message[110] ^ CRC_i_Message[111] ^ CRC_i_Message[113] ^ CRC_i_Message[117] ^ CRC_i_Message[120] ^ CRC_i_Message[125] ^ CRC_i_Message[126]);
			CRC_o_CRC[30] = ~(temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 40] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 90] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[105] ^ CRC_i_Message[106] ^ CRC_i_Message[108] ^ CRC_i_Message[109] ^ CRC_i_Message[110] ^ CRC_i_Message[112] ^ CRC_i_Message[116] ^ CRC_i_Message[119] ^ CRC_i_Message[124] ^ CRC_i_Message[125]);
			CRC_o_CRC[29] = ~(temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  8] ^ temp_seed[  9] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 21] ^ temp_seed[ 23] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 39] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 54] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 89] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 99] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[105] ^ CRC_i_Message[107] ^ CRC_i_Message[108] ^ CRC_i_Message[109] ^ CRC_i_Message[117] ^ CRC_i_Message[121] ^ CRC_i_Message[123] ^ CRC_i_Message[124] ^ CRC_i_Message[127]);
			CRC_o_CRC[28] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  9] ^ temp_seed[ 10] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 22] ^ temp_seed[ 24] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  7] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 38] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 53] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 88] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 98] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[106] ^ CRC_i_Message[107] ^ CRC_i_Message[108] ^ CRC_i_Message[116] ^ CRC_i_Message[120] ^ CRC_i_Message[122] ^ CRC_i_Message[123] ^ CRC_i_Message[126]);
			CRC_o_CRC[27] = ~(temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[ 10] ^ temp_seed[ 11] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 23] ^ temp_seed[ 25] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  6] ^ CRC_i_Message[  8] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 21] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 37] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 52] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 59] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 87] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[105] ^ CRC_i_Message[106] ^ CRC_i_Message[107] ^ CRC_i_Message[115] ^ CRC_i_Message[119] ^ CRC_i_Message[121] ^ CRC_i_Message[122] ^ CRC_i_Message[125]);
			CRC_o_CRC[26] = ~(temp_seed[  0] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  5] ^ temp_seed[  7] ^ temp_seed[ 11] ^ temp_seed[ 12] ^ temp_seed[ 14] ^ temp_seed[ 15] ^ temp_seed[ 17] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 24] ^ temp_seed[ 26] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  5] ^ CRC_i_Message[  7] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 20] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 36] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 51] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 58] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 72] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 77] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 86] ^ CRC_i_Message[ 93] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[102] ^ CRC_i_Message[104] ^ CRC_i_Message[105] ^ CRC_i_Message[106] ^ CRC_i_Message[114] ^ CRC_i_Message[118] ^ CRC_i_Message[120] ^ CRC_i_Message[121] ^ CRC_i_Message[124]);
			CRC_o_CRC[25] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  3] ^ temp_seed[  5] ^ temp_seed[  6] ^ temp_seed[  8] ^ temp_seed[ 12] ^ temp_seed[ 13] ^ temp_seed[ 15] ^ temp_seed[ 16] ^ temp_seed[ 18] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 25] ^ temp_seed[ 27] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  4] ^ CRC_i_Message[  6] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 13] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 16] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 19] ^ CRC_i_Message[ 23] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 26] ^ CRC_i_Message[ 28] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 35] ^ CRC_i_Message[ 42] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 48] ^ CRC_i_Message[ 50] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 57] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 64] ^ CRC_i_Message[ 66] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 69] ^ CRC_i_Message[ 71] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 76] ^ CRC_i_Message[ 79] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 82] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 85] ^ CRC_i_Message[ 92] ^ CRC_i_Message[ 95] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[101] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[105] ^ CRC_i_Message[113] ^ CRC_i_Message[117] ^ CRC_i_Message[119] ^ CRC_i_Message[120] ^ CRC_i_Message[123]);
			CRC_o_CRC[24] = ~(temp_seed[  0] ^ temp_seed[  1] ^ temp_seed[  2] ^ temp_seed[  4] ^ temp_seed[  6] ^ temp_seed[  7] ^ temp_seed[  9] ^ temp_seed[ 13] ^ temp_seed[ 14] ^ temp_seed[ 16] ^ temp_seed[ 17] ^ temp_seed[ 19] ^ temp_seed[ 20] ^ temp_seed[ 21] ^ temp_seed[ 22] ^ temp_seed[ 26] ^ temp_seed[ 28] ^ temp_seed[ 29] ^ temp_seed[ 30] ^ temp_seed[ 31] ^ CRC_i_Message[  0] ^ CRC_i_Message[  1] ^ CRC_i_Message[  2] ^ CRC_i_Message[  3] ^ CRC_i_Message[  5] ^ CRC_i_Message[  9] ^ CRC_i_Message[ 10] ^ CRC_i_Message[ 11] ^ CRC_i_Message[ 12] ^ CRC_i_Message[ 14] ^ CRC_i_Message[ 15] ^ CRC_i_Message[ 17] ^ CRC_i_Message[ 18] ^ CRC_i_Message[ 22] ^ CRC_i_Message[ 24] ^ CRC_i_Message[ 25] ^ CRC_i_Message[ 27] ^ CRC_i_Message[ 29] ^ CRC_i_Message[ 30] ^ CRC_i_Message[ 31] ^ CRC_i_Message[ 32] ^ CRC_i_Message[ 33] ^ CRC_i_Message[ 34] ^ CRC_i_Message[ 41] ^ CRC_i_Message[ 43] ^ CRC_i_Message[ 44] ^ CRC_i_Message[ 45] ^ CRC_i_Message[ 46] ^ CRC_i_Message[ 47] ^ CRC_i_Message[ 49] ^ CRC_i_Message[ 55] ^ CRC_i_Message[ 56] ^ CRC_i_Message[ 60] ^ CRC_i_Message[ 61] ^ CRC_i_Message[ 62] ^ CRC_i_Message[ 63] ^ CRC_i_Message[ 65] ^ CRC_i_Message[ 67] ^ CRC_i_Message[ 68] ^ CRC_i_Message[ 70] ^ CRC_i_Message[ 73] ^ CRC_i_Message[ 74] ^ CRC_i_Message[ 75] ^ CRC_i_Message[ 78] ^ CRC_i_Message[ 80] ^ CRC_i_Message[ 81] ^ CRC_i_Message[ 83] ^ CRC_i_Message[ 84] ^ CRC_i_Message[ 91] ^ CRC_i_Message[ 94] ^ CRC_i_Message[ 96] ^ CRC_i_Message[ 97] ^ CRC_i_Message[ 98] ^ CRC_i_Message[ 99] ^ CRC_i_Message[100] ^ CRC_i_Message[102] ^ CRC_i_Message[103] ^ CRC_i_Message[104] ^ CRC_i_Message[112] ^ CRC_i_Message[116] ^ CRC_i_Message[118] ^ CRC_i_Message[119] ^ CRC_i_Message[122]);
		end
		// Data Length 160 bits (5DW)
		else if (CRC_i_Length == 'd5) begin
			CRC_o_CRC[ 7] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[159] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 6] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[135] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[65] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[21] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 5] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[115] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 4] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[114] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[83] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3]);
			CRC_o_CRC[ 3] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[144] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 2] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[146] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 1] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[145] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[134] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 0] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[72] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[3] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[15] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[142] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[14] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[141] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[13] = ~(temp_seed[2] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[12] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[46] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3]);
			CRC_o_CRC[11] = ~(temp_seed[0] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[18] ^ CRC_i_Message[14] ^ CRC_i_Message[10] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[10] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[134] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[17] ^ CRC_i_Message[13] ^ CRC_i_Message[9] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 9] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[133] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[16] ^ CRC_i_Message[12] ^ CRC_i_Message[8] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 8] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[15] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[23] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[159] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[28] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[22] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[158] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[21] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[157] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[20] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[156] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[19] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[155] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[18] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[154] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[17] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[80] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[16] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[89] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[30] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[29] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[28] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[149] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[3]);
			CRC_o_CRC[28] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[148] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[27] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[147] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[26] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[156] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[25] = ~(temp_seed[2] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[31] ^ CRC_i_Message[155] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[0]);
			CRC_o_CRC[24] = ~(temp_seed[3] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2]);
		end	
        // Data Length 192 bits	(6DW)
		else if (CRC_i_Length == 'd6) begin
			CRC_o_CRC[ 7] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[6] 	^ temp_seed[7]  ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[191] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[175] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 6] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[6] 	^ temp_seed[8]  ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[167] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[97] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[53] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[18] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 5] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] 	^ temp_seed[6]  ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[147] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2]);
			CRC_o_CRC[ 4] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] 	^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[146] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[8] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 3] = ~(temp_seed[3] ^ temp_seed[7] ^ temp_seed[8] 	^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[176] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[28] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 2] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[4] 	^ temp_seed[6]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[178] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4]);
			CRC_o_CRC[ 1] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] 	^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[177] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[166] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3]);
			CRC_o_CRC[ 0] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] 	^ temp_seed[7]  ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[104] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[15] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] 	^ temp_seed[3]  ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[174] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5]);
			CRC_o_CRC[14] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] 	^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[173] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4]);
			CRC_o_CRC[13] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] 	^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[182] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[172] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[12] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[5] 	^ temp_seed[7]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[30] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[171] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[97] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[78] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[1]);
			CRC_o_CRC[11] = ~(temp_seed[2] ^ temp_seed[5] ^ temp_seed[7] 	^ temp_seed[8]  ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[164] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[86] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[46] ^ CRC_i_Message[42] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[10] = ~(temp_seed[3] ^ temp_seed[6] ^ temp_seed[8] 	^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[169] ^ CRC_i_Message[166] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[49] ^ CRC_i_Message[45] ^ CRC_i_Message[41] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[28] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 9] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[7] 	^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[168] ^ CRC_i_Message[165] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[44] ^ CRC_i_Message[40] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 8] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5] 	^ temp_seed[8]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[164] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[83] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[47] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[23] = ~(temp_seed[0] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[191] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[183] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[22] = ~(temp_seed[1] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[190] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[21] = ~(temp_seed[2] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[31] ^ CRC_i_Message[189] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[0]);
			CRC_o_CRC[20] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[188] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[28] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[19] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4]  ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[187] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[20] ^ CRC_i_Message[17] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[18] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2]  ^ temp_seed[5]  ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[186] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[178] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[17] = ~(temp_seed[3] ^ temp_seed[7] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ CRC_i_Message[191] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[112] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[28] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2]);
			CRC_o_CRC[16] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2]  ^ temp_seed[4]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[31] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[14] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2]  ^ temp_seed[3]  ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[3]);
			CRC_o_CRC[30] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3]  ^ temp_seed[4]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[2]);
			CRC_o_CRC[29] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3]  ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[31] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[181] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[0]);
			CRC_o_CRC[28] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[180] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[27] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[189] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[179] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[26] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[6]  ^ temp_seed[7]  ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[188] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[178] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[25] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[7]  ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[187] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[177] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[24] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5]  ^ temp_seed[6]  ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[186] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
		end	
        // Data Length 224 bits	(7DW)
		else if (CRC_i_Length == 'd7) begin
			CRC_o_CRC[ 7] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^CRC_i_Message[223] ^ CRC_i_Message[217] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[211] ^ CRC_i_Message[207] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[186] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[7]);
			CRC_o_CRC[ 6] = ~(temp_seed[3] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9]  ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[199] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[129] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[103] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[85] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6]);
			CRC_o_CRC[ 5] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[179] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[121] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[41] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5]);
			CRC_o_CRC[ 4] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[178] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[40] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4]);
			CRC_o_CRC[ 3] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^CRC_i_Message[223] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[217] ^ CRC_i_Message[215] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[208] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[60] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3]);
			CRC_o_CRC[ 2] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[213] ^ CRC_i_Message[210] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[199] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[ 1] = ~(temp_seed[1] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[212] ^ CRC_i_Message[209] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[198] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[119] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 0] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5] ^ temp_seed[7]  ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[223] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[136] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[15] = ~(temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[206] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[195] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[14] = ~(temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[205] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[194] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[17] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[13] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[223] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[214] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[204] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[19] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[12] = ~(temp_seed[3] ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[214] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[203] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[110] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[63] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[33] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[11] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[214] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[202] ^ CRC_i_Message[199] ^ CRC_i_Message[196] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[82] ^ CRC_i_Message[78] ^ CRC_i_Message[74] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[10] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[213] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[201] ^ CRC_i_Message[198] ^ CRC_i_Message[195] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[81] ^ CRC_i_Message[77] ^ CRC_i_Message[73] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 9] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[212] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[200] ^ CRC_i_Message[197] ^ CRC_i_Message[194] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[116] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[76] ^ CRC_i_Message[72] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 8] = ~(temp_seed[1] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[211] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[199] ^ CRC_i_Message[196] ^ CRC_i_Message[193] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[115] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[79] ^ CRC_i_Message[75] ^ CRC_i_Message[71] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[23] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[8]  ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[223] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[215] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[206] ^ CRC_i_Message[204] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[172] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[22] = ~(temp_seed[2] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9]  ^ temp_seed[11] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[222] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[214] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[205] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[171] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[21] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[9]  ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[221] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[213] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[204] ^ CRC_i_Message[202] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[170] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[28] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[20] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[7]  ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[220] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[212] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[169] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[19] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[8]  ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[219] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[211] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[202] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[168] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[18] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[6] ^ temp_seed[9]  ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[218] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[210] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[17] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[30] ^ CRC_i_Message[223] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[171] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[144] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[60] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[1]);
			CRC_o_CRC[16] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[31] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[217] ^ CRC_i_Message[214] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[36] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[216] ^ CRC_i_Message[213] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3]);
			CRC_o_CRC[30] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[215] ^ CRC_i_Message[212] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[34] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[29] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[223] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[217] ^ CRC_i_Message[213] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[192] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[28] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4]  ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[222] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[212] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[191] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[27] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[221] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[215] ^ CRC_i_Message[211] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[190] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[26] = ~(temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[6]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[220] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[214] ^ CRC_i_Message[210] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[189] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[25] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[30] ^ CRC_i_Message[219] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[209] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[1]);
			CRC_o_CRC[24] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[5]  ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[31] ^ CRC_i_Message[218] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[208] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[0]);
		end	
        // Data Length 256 bits	(8DW)
		else if (CRC_i_Length == 'd8) begin
			CRC_o_CRC[ 7] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[19] ^ temp_seed[24] ^ temp_seed[28] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[249] ^ CRC_i_Message[246] ^ CRC_i_Message[245] ^ CRC_i_Message[243] ^ CRC_i_Message[239] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[225] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[221] ^ CRC_i_Message[218] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[12] ^ CRC_i_Message[7] ^ CRC_i_Message[3] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 6] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[246] ^ CRC_i_Message[244] ^ CRC_i_Message[243] ^ CRC_i_Message[242] ^ CRC_i_Message[239] ^ CRC_i_Message[238] ^ CRC_i_Message[231] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[202] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[186] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[161] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[135] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[117] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[82] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 5] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[246] ^ CRC_i_Message[242] ^ CRC_i_Message[241] ^ CRC_i_Message[239] ^ CRC_i_Message[238] ^ CRC_i_Message[237] ^ CRC_i_Message[231] ^ CRC_i_Message[229] ^ CRC_i_Message[225] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[211] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[153] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[109] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[73] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 4] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[246] ^ CRC_i_Message[245] ^ CRC_i_Message[241] ^ CRC_i_Message[240] ^ CRC_i_Message[238] ^ CRC_i_Message[237] ^ CRC_i_Message[236] ^ CRC_i_Message[230] ^ CRC_i_Message[228] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[210] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[190] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[179] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[152] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[72] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 3] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[30] ^ CRC_i_Message[255] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[249] ^ CRC_i_Message[247] ^ CRC_i_Message[244] ^ CRC_i_Message[243] ^ CRC_i_Message[240] ^ CRC_i_Message[237] ^ CRC_i_Message[236] ^ CRC_i_Message[235] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[226] ^ CRC_i_Message[225] ^ CRC_i_Message[224] ^ CRC_i_Message[222] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[92] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 2] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[27] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[245] ^ CRC_i_Message[242] ^ CRC_i_Message[236] ^ CRC_i_Message[235] ^ CRC_i_Message[234] ^ CRC_i_Message[231] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[63] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[4]);
			CRC_o_CRC[ 1] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[28] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[244] ^ CRC_i_Message[241] ^ CRC_i_Message[235] ^ CRC_i_Message[234] ^ CRC_i_Message[233] ^ CRC_i_Message[230] ^ CRC_i_Message[226] ^ CRC_i_Message[225] ^ CRC_i_Message[217] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[62] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[3]);
			CRC_o_CRC[ 0] = ~(temp_seed[0] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[250] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[245] ^ CRC_i_Message[240] ^ CRC_i_Message[239] ^ CRC_i_Message[234] ^ CRC_i_Message[233] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[223] ^ CRC_i_Message[221] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[168] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[18] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[15] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[247] ^ CRC_i_Message[245] ^ CRC_i_Message[244] ^ CRC_i_Message[243] ^ CRC_i_Message[238] ^ CRC_i_Message[233] ^ CRC_i_Message[232] ^ CRC_i_Message[227] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[14] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[246] ^ CRC_i_Message[244] ^ CRC_i_Message[243] ^ CRC_i_Message[242] ^ CRC_i_Message[237] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[226] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[200] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[81] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[12] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[13] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ CRC_i_Message[255] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[250] ^ CRC_i_Message[246] ^ CRC_i_Message[242] ^ CRC_i_Message[241] ^ CRC_i_Message[239] ^ CRC_i_Message[236] ^ CRC_i_Message[229] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[205] ^ CRC_i_Message[203] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[189] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[172] ^ CRC_i_Message[169] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[82] ^ CRC_i_Message[80] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[51] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5]);
			CRC_o_CRC[12] = ~(temp_seed[1] ^ temp_seed[4] ^ temp_seed[10] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[246] ^ CRC_i_Message[243] ^ CRC_i_Message[241] ^ CRC_i_Message[240] ^ CRC_i_Message[239] ^ CRC_i_Message[238] ^ CRC_i_Message[235] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[224] ^ CRC_i_Message[222] ^ CRC_i_Message[219] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[161] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[142] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[121] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[95] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[81] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[65] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[21] ^ CRC_i_Message[19] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[0]);
			CRC_o_CRC[11] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[249] ^ CRC_i_Message[246] ^ CRC_i_Message[243] ^ CRC_i_Message[242] ^ CRC_i_Message[240] ^ CRC_i_Message[238] ^ CRC_i_Message[237] ^ CRC_i_Message[234] ^ CRC_i_Message[231] ^ CRC_i_Message[228] ^ CRC_i_Message[225] ^ CRC_i_Message[224] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[114] ^ CRC_i_Message[110] ^ CRC_i_Message[106] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[80] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[10] = ~(temp_seed[4] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[250] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[245] ^ CRC_i_Message[242] ^ CRC_i_Message[241] ^ CRC_i_Message[239] ^ CRC_i_Message[237] ^ CRC_i_Message[236] ^ CRC_i_Message[233] ^ CRC_i_Message[230] ^ CRC_i_Message[227] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[149] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[113] ^ CRC_i_Message[109] ^ CRC_i_Message[105] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[92] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[79] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[ 9] = ~(temp_seed[0] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[244] ^ CRC_i_Message[241] ^ CRC_i_Message[240] ^ CRC_i_Message[238] ^ CRC_i_Message[236] ^ CRC_i_Message[235] ^ CRC_i_Message[232] ^ CRC_i_Message[229] ^ CRC_i_Message[226] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[190] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[148] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[112] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[91] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[78] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[63] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[ 8] = ~(temp_seed[1] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[30] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[246] ^ CRC_i_Message[243] ^ CRC_i_Message[240] ^ CRC_i_Message[239] ^ CRC_i_Message[237] ^ CRC_i_Message[235] ^ CRC_i_Message[234] ^ CRC_i_Message[231] ^ CRC_i_Message[228] ^ CRC_i_Message[225] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[189] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[111] ^ CRC_i_Message[107] ^ CRC_i_Message[103] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[90] ^ CRC_i_Message[87] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[77] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[42] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[1]);
			
			CRC_o_CRC[23] = ~(temp_seed[3] ^ temp_seed[4] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ CRC_i_Message[255] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[247] ^ CRC_i_Message[243] ^ CRC_i_Message[242] ^ CRC_i_Message[238] ^ CRC_i_Message[236] ^ CRC_i_Message[234] ^ CRC_i_Message[233] ^ CRC_i_Message[231] ^ CRC_i_Message[229] ^ CRC_i_Message[226] ^ CRC_i_Message[225] ^ CRC_i_Message[223] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[204] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[189] ^ CRC_i_Message[187] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[88] ^ CRC_i_Message[85] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[76] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[53] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5]);
			CRC_o_CRC[22] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ CRC_i_Message[254] ^ CRC_i_Message[250] ^ CRC_i_Message[249] ^ CRC_i_Message[246] ^ CRC_i_Message[242] ^ CRC_i_Message[241] ^ CRC_i_Message[237] ^ CRC_i_Message[235] ^ CRC_i_Message[233] ^ CRC_i_Message[232] ^ CRC_i_Message[230] ^ CRC_i_Message[228] ^ CRC_i_Message[225] ^ CRC_i_Message[224] ^ CRC_i_Message[222] ^ CRC_i_Message[219] ^ CRC_i_Message[217] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[203] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[188] ^ CRC_i_Message[186] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[94] ^ CRC_i_Message[87] ^ CRC_i_Message[84] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4]);
			CRC_o_CRC[21] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[28] ^ CRC_i_Message[253] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[245] ^ CRC_i_Message[241] ^ CRC_i_Message[240] ^ CRC_i_Message[236] ^ CRC_i_Message[234] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[229] ^ CRC_i_Message[227] ^ CRC_i_Message[224] ^ CRC_i_Message[223] ^ CRC_i_Message[221] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[202] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[187] ^ CRC_i_Message[185] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[93] ^ CRC_i_Message[86] ^ CRC_i_Message[83] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[3]);
			CRC_o_CRC[20] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[6] ^ temp_seed[7] ^ temp_seed[9] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[29] ^ CRC_i_Message[252] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[244] ^ CRC_i_Message[240] ^ CRC_i_Message[239] ^ CRC_i_Message[235] ^ CRC_i_Message[233] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[228] ^ CRC_i_Message[226] ^ CRC_i_Message[223] ^ CRC_i_Message[222] ^ CRC_i_Message[220] ^ CRC_i_Message[217] ^ CRC_i_Message[215] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[201] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[186] ^ CRC_i_Message[184] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[128] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[121] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[92] ^ CRC_i_Message[85] ^ CRC_i_Message[82] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[56] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[25] ^ CRC_i_Message[24] ^ CRC_i_Message[22] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[2]);
			CRC_o_CRC[19] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[7] ^ temp_seed[8] ^ temp_seed[10] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[30] ^ CRC_i_Message[251] ^ CRC_i_Message[247] ^ CRC_i_Message[246] ^ CRC_i_Message[243] ^ CRC_i_Message[239] ^ CRC_i_Message[238] ^ CRC_i_Message[234] ^ CRC_i_Message[232] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[227] ^ CRC_i_Message[225] ^ CRC_i_Message[222] ^ CRC_i_Message[221] ^ CRC_i_Message[219] ^ CRC_i_Message[216] ^ CRC_i_Message[214] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[200] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[185] ^ CRC_i_Message[183] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[127] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[120] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[113] ^ CRC_i_Message[111] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[91] ^ CRC_i_Message[84] ^ CRC_i_Message[81] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[58] ^ CRC_i_Message[55] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[24] ^ CRC_i_Message[23] ^ CRC_i_Message[21] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[1]);
			CRC_o_CRC[18] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[8] ^ temp_seed[9] ^ temp_seed[11] ^ temp_seed[12] ^ temp_seed[13] ^ temp_seed[14] ^ temp_seed[18] ^ temp_seed[19] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[250] ^ CRC_i_Message[246] ^ CRC_i_Message[245] ^ CRC_i_Message[242] ^ CRC_i_Message[238] ^ CRC_i_Message[237] ^ CRC_i_Message[233] ^ CRC_i_Message[231] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[226] ^ CRC_i_Message[224] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[218] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[206] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[199] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[184] ^ CRC_i_Message[182] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[156] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[126] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[119] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[90] ^ CRC_i_Message[83] ^ CRC_i_Message[80] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[57] ^ CRC_i_Message[54] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[23] ^ CRC_i_Message[22] ^ CRC_i_Message[20] ^ CRC_i_Message[19] ^ CRC_i_Message[18] ^ CRC_i_Message[17] ^ CRC_i_Message[13] ^ CRC_i_Message[12] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			CRC_o_CRC[17] = ~(temp_seed[1] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[14] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[21] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ CRC_i_Message[255] ^ CRC_i_Message[246] ^ CRC_i_Message[244] ^ CRC_i_Message[243] ^ CRC_i_Message[241] ^ CRC_i_Message[239] ^ CRC_i_Message[237] ^ CRC_i_Message[236] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[226] ^ CRC_i_Message[224] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[203] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[176] ^ CRC_i_Message[173] ^ CRC_i_Message[170] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[109] ^ CRC_i_Message[108] ^ CRC_i_Message[105] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[92] ^ CRC_i_Message[88] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[83] ^ CRC_i_Message[82] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[45] ^ CRC_i_Message[44] ^ CRC_i_Message[43] ^ CRC_i_Message[42] ^ CRC_i_Message[41] ^ CRC_i_Message[40] ^ CRC_i_Message[39] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[33] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[17] ^ CRC_i_Message[16] ^ CRC_i_Message[11] ^ CRC_i_Message[10] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[2]);
			CRC_o_CRC[16] = ~(temp_seed[0] ^ temp_seed[3] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[15] ^ temp_seed[16] ^ temp_seed[19] ^ temp_seed[21] ^ temp_seed[22] ^ temp_seed[24] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[30] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[254] ^ CRC_i_Message[249] ^ CRC_i_Message[246] ^ CRC_i_Message[242] ^ CRC_i_Message[240] ^ CRC_i_Message[239] ^ CRC_i_Message[238] ^ CRC_i_Message[236] ^ CRC_i_Message[235] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[226] ^ CRC_i_Message[224] ^ CRC_i_Message[221] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[213] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[190] ^ CRC_i_Message[186] ^ CRC_i_Message[183] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[162] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[120] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[108] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[82] ^ CRC_i_Message[81] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[68] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[54] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[28] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[16] ^ CRC_i_Message[15] ^ CRC_i_Message[12] ^ CRC_i_Message[10] ^ CRC_i_Message[9] ^ CRC_i_Message[7] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[1] ^ CRC_i_Message[0]);
			
			CRC_o_CRC[31] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[4] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[16] ^ temp_seed[17] ^ temp_seed[20] ^ temp_seed[22] ^ temp_seed[23] ^ temp_seed[25] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[31] ^ CRC_i_Message[254] ^ CRC_i_Message[253] ^ CRC_i_Message[248] ^ CRC_i_Message[245] ^ CRC_i_Message[241] ^ CRC_i_Message[239] ^ CRC_i_Message[238] ^ CRC_i_Message[237] ^ CRC_i_Message[235] ^ CRC_i_Message[234] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[225] ^ CRC_i_Message[223] ^ CRC_i_Message[220] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[212] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[189] ^ CRC_i_Message[185] ^ CRC_i_Message[182] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[161] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[139] ^ CRC_i_Message[137] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[130] ^ CRC_i_Message[128] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[119] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[107] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[99] ^ CRC_i_Message[97] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[81] ^ CRC_i_Message[80] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[67] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[53] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[39] ^ CRC_i_Message[37] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[27] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[15] ^ CRC_i_Message[14] ^ CRC_i_Message[11] ^ CRC_i_Message[9] ^ CRC_i_Message[8] ^ CRC_i_Message[6] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[0]);
			CRC_o_CRC[30] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[5] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[17] ^ temp_seed[18] ^ temp_seed[21] ^ temp_seed[23] ^ temp_seed[24] ^ temp_seed[26] ^ temp_seed[27] ^ temp_seed[28] ^ CRC_i_Message[253] ^ CRC_i_Message[252] ^ CRC_i_Message[247] ^ CRC_i_Message[244] ^ CRC_i_Message[240] ^ CRC_i_Message[238] ^ CRC_i_Message[237] ^ CRC_i_Message[236] ^ CRC_i_Message[234] ^ CRC_i_Message[233] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[224] ^ CRC_i_Message[222] ^ CRC_i_Message[219] ^ CRC_i_Message[218] ^ CRC_i_Message[217] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[211] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[188] ^ CRC_i_Message[184] ^ CRC_i_Message[181] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[168] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[118] ^ CRC_i_Message[112] ^ CRC_i_Message[111] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[98] ^ CRC_i_Message[96] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[80] ^ CRC_i_Message[79] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[72] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[66] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[52] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[38] ^ CRC_i_Message[36] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[26] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[14] ^ CRC_i_Message[13] ^ CRC_i_Message[10] ^ CRC_i_Message[8] ^ CRC_i_Message[7] ^ CRC_i_Message[5] ^ CRC_i_Message[4] ^ CRC_i_Message[3]);
			CRC_o_CRC[29] = ~(temp_seed[0] ^ temp_seed[4] ^ temp_seed[7] ^ temp_seed[13] ^ temp_seed[18] ^ temp_seed[22] ^ temp_seed[25] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[255] ^ CRC_i_Message[252] ^ CRC_i_Message[251] ^ CRC_i_Message[249] ^ CRC_i_Message[245] ^ CRC_i_Message[237] ^ CRC_i_Message[236] ^ CRC_i_Message[235] ^ CRC_i_Message[233] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[227] ^ CRC_i_Message[224] ^ CRC_i_Message[217] ^ CRC_i_Message[216] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[211] ^ CRC_i_Message[208] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[203] ^ CRC_i_Message[201] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[182] ^ CRC_i_Message[180] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[174] ^ CRC_i_Message[167] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[151] ^ CRC_i_Message[150] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[138] ^ CRC_i_Message[136] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[129] ^ CRC_i_Message[127] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[118] ^ CRC_i_Message[117] ^ CRC_i_Message[112] ^ CRC_i_Message[110] ^ CRC_i_Message[106] ^ CRC_i_Message[105] ^ CRC_i_Message[103] ^ CRC_i_Message[100] ^ CRC_i_Message[99] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[79] ^ CRC_i_Message[78] ^ CRC_i_Message[75] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[37] ^ CRC_i_Message[35] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[27] ^ CRC_i_Message[24] ^ CRC_i_Message[18] ^ CRC_i_Message[13] ^ CRC_i_Message[9] ^ CRC_i_Message[6] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[28] = ~(temp_seed[1] ^ temp_seed[5] ^ temp_seed[8] ^ temp_seed[14] ^ temp_seed[19] ^ temp_seed[23] ^ temp_seed[26] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[254] ^ CRC_i_Message[251] ^ CRC_i_Message[250] ^ CRC_i_Message[248] ^ CRC_i_Message[244] ^ CRC_i_Message[236] ^ CRC_i_Message[235] ^ CRC_i_Message[234] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[226] ^ CRC_i_Message[223] ^ CRC_i_Message[216] ^ CRC_i_Message[215] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[210] ^ CRC_i_Message[207] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[202] ^ CRC_i_Message[200] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[188] ^ CRC_i_Message[187] ^ CRC_i_Message[181] ^ CRC_i_Message[179] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[173] ^ CRC_i_Message[166] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[150] ^ CRC_i_Message[149] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[137] ^ CRC_i_Message[135] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[128] ^ CRC_i_Message[126] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[117] ^ CRC_i_Message[116] ^ CRC_i_Message[111] ^ CRC_i_Message[109] ^ CRC_i_Message[105] ^ CRC_i_Message[104] ^ CRC_i_Message[102] ^ CRC_i_Message[99] ^ CRC_i_Message[98] ^ CRC_i_Message[94] ^ CRC_i_Message[93] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[78] ^ CRC_i_Message[77] ^ CRC_i_Message[74] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[53] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[36] ^ CRC_i_Message[34] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[26] ^ CRC_i_Message[23] ^ CRC_i_Message[17] ^ CRC_i_Message[12] ^ CRC_i_Message[8] ^ CRC_i_Message[5] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[27] = ~(temp_seed[0] ^ temp_seed[2] ^ temp_seed[6] ^ temp_seed[9] ^ temp_seed[15] ^ temp_seed[20] ^ temp_seed[24] ^ temp_seed[27] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[253] ^ CRC_i_Message[250] ^ CRC_i_Message[249] ^ CRC_i_Message[247] ^ CRC_i_Message[243] ^ CRC_i_Message[235] ^ CRC_i_Message[234] ^ CRC_i_Message[233] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[225] ^ CRC_i_Message[222] ^ CRC_i_Message[215] ^ CRC_i_Message[214] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[206] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[201] ^ CRC_i_Message[199] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[187] ^ CRC_i_Message[186] ^ CRC_i_Message[180] ^ CRC_i_Message[178] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[172] ^ CRC_i_Message[165] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[149] ^ CRC_i_Message[148] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[136] ^ CRC_i_Message[134] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[127] ^ CRC_i_Message[125] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[116] ^ CRC_i_Message[115] ^ CRC_i_Message[110] ^ CRC_i_Message[108] ^ CRC_i_Message[104] ^ CRC_i_Message[103] ^ CRC_i_Message[101] ^ CRC_i_Message[98] ^ CRC_i_Message[97] ^ CRC_i_Message[93] ^ CRC_i_Message[92] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[77] ^ CRC_i_Message[76] ^ CRC_i_Message[73] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[62] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[52] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[35] ^ CRC_i_Message[33] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[29] ^ CRC_i_Message[25] ^ CRC_i_Message[22] ^ CRC_i_Message[16] ^ CRC_i_Message[11] ^ CRC_i_Message[7] ^ CRC_i_Message[4] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[26] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[3] ^ temp_seed[7] ^ temp_seed[10] ^ temp_seed[16] ^ temp_seed[21] ^ temp_seed[25] ^ temp_seed[28] ^ temp_seed[30] ^ CRC_i_Message[252] ^ CRC_i_Message[249] ^ CRC_i_Message[248] ^ CRC_i_Message[246] ^ CRC_i_Message[242] ^ CRC_i_Message[234] ^ CRC_i_Message[233] ^ CRC_i_Message[232] ^ CRC_i_Message[230] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[224] ^ CRC_i_Message[221] ^ CRC_i_Message[214] ^ CRC_i_Message[213] ^ CRC_i_Message[211] ^ CRC_i_Message[210] ^ CRC_i_Message[208] ^ CRC_i_Message[205] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[200] ^ CRC_i_Message[198] ^ CRC_i_Message[197] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[186] ^ CRC_i_Message[185] ^ CRC_i_Message[179] ^ CRC_i_Message[177] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[171] ^ CRC_i_Message[164] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[154] ^ CRC_i_Message[152] ^ CRC_i_Message[148] ^ CRC_i_Message[147] ^ CRC_i_Message[145] ^ CRC_i_Message[144] ^ CRC_i_Message[142] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[135] ^ CRC_i_Message[133] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[126] ^ CRC_i_Message[124] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[115] ^ CRC_i_Message[114] ^ CRC_i_Message[109] ^ CRC_i_Message[107] ^ CRC_i_Message[103] ^ CRC_i_Message[102] ^ CRC_i_Message[100] ^ CRC_i_Message[97] ^ CRC_i_Message[96] ^ CRC_i_Message[92] ^ CRC_i_Message[91] ^ CRC_i_Message[89] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[76] ^ CRC_i_Message[75] ^ CRC_i_Message[72] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[61] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[57] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[51] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[34] ^ CRC_i_Message[32] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[28] ^ CRC_i_Message[24] ^ CRC_i_Message[21] ^ CRC_i_Message[15] ^ CRC_i_Message[10] ^ CRC_i_Message[6] ^ CRC_i_Message[3] ^ CRC_i_Message[1]);
			CRC_o_CRC[25] = ~(temp_seed[0] ^ temp_seed[1] ^ temp_seed[2] ^ temp_seed[4] ^ temp_seed[8] ^ temp_seed[11] ^ temp_seed[17] ^ temp_seed[22] ^ temp_seed[26] ^ temp_seed[29] ^ temp_seed[31] ^ CRC_i_Message[251] ^ CRC_i_Message[248] ^ CRC_i_Message[247] ^ CRC_i_Message[245] ^ CRC_i_Message[241] ^ CRC_i_Message[233] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[229] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[225] ^ CRC_i_Message[223] ^ CRC_i_Message[220] ^ CRC_i_Message[213] ^ CRC_i_Message[212] ^ CRC_i_Message[210] ^ CRC_i_Message[209] ^ CRC_i_Message[207] ^ CRC_i_Message[204] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[199] ^ CRC_i_Message[197] ^ CRC_i_Message[196] ^ CRC_i_Message[194] ^ CRC_i_Message[192] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[185] ^ CRC_i_Message[184] ^ CRC_i_Message[178] ^ CRC_i_Message[176] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[170] ^ CRC_i_Message[163] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[156] ^ CRC_i_Message[154] ^ CRC_i_Message[153] ^ CRC_i_Message[151] ^ CRC_i_Message[147] ^ CRC_i_Message[146] ^ CRC_i_Message[144] ^ CRC_i_Message[143] ^ CRC_i_Message[141] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[134] ^ CRC_i_Message[132] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[125] ^ CRC_i_Message[123] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[114] ^ CRC_i_Message[113] ^ CRC_i_Message[108] ^ CRC_i_Message[106] ^ CRC_i_Message[102] ^ CRC_i_Message[101] ^ CRC_i_Message[99] ^ CRC_i_Message[96] ^ CRC_i_Message[95] ^ CRC_i_Message[91] ^ CRC_i_Message[90] ^ CRC_i_Message[88] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[75] ^ CRC_i_Message[74] ^ CRC_i_Message[71] ^ CRC_i_Message[69] ^ CRC_i_Message[67] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[60] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[56] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[50] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[45] ^ CRC_i_Message[43] ^ CRC_i_Message[41] ^ CRC_i_Message[33] ^ CRC_i_Message[31] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[27] ^ CRC_i_Message[23] ^ CRC_i_Message[20] ^ CRC_i_Message[14] ^ CRC_i_Message[9] ^ CRC_i_Message[5] ^ CRC_i_Message[2] ^ CRC_i_Message[0]);
			CRC_o_CRC[24] = ~(temp_seed[1] ^ temp_seed[2] ^ temp_seed[3] ^ temp_seed[5] ^ temp_seed[9] ^ temp_seed[12] ^ temp_seed[18] ^ temp_seed[23] ^ temp_seed[27] ^ temp_seed[30] ^ CRC_i_Message[250] ^ CRC_i_Message[247] ^ CRC_i_Message[246] ^ CRC_i_Message[244] ^ CRC_i_Message[240] ^ CRC_i_Message[232] ^ CRC_i_Message[231] ^ CRC_i_Message[230] ^ CRC_i_Message[228] ^ CRC_i_Message[227] ^ CRC_i_Message[226] ^ CRC_i_Message[225] ^ CRC_i_Message[224] ^ CRC_i_Message[222] ^ CRC_i_Message[219] ^ CRC_i_Message[212] ^ CRC_i_Message[211] ^ CRC_i_Message[209] ^ CRC_i_Message[208] ^ CRC_i_Message[206] ^ CRC_i_Message[203] ^ CRC_i_Message[202] ^ CRC_i_Message[201] ^ CRC_i_Message[198] ^ CRC_i_Message[196] ^ CRC_i_Message[195] ^ CRC_i_Message[193] ^ CRC_i_Message[191] ^ CRC_i_Message[190] ^ CRC_i_Message[189] ^ CRC_i_Message[188] ^ CRC_i_Message[184] ^ CRC_i_Message[183] ^ CRC_i_Message[177] ^ CRC_i_Message[175] ^ CRC_i_Message[174] ^ CRC_i_Message[173] ^ CRC_i_Message[172] ^ CRC_i_Message[171] ^ CRC_i_Message[169] ^ CRC_i_Message[162] ^ CRC_i_Message[161] ^ CRC_i_Message[160] ^ CRC_i_Message[159] ^ CRC_i_Message[158] ^ CRC_i_Message[157] ^ CRC_i_Message[155] ^ CRC_i_Message[153] ^ CRC_i_Message[152] ^ CRC_i_Message[150] ^ CRC_i_Message[146] ^ CRC_i_Message[145] ^ CRC_i_Message[143] ^ CRC_i_Message[142] ^ CRC_i_Message[140] ^ CRC_i_Message[139] ^ CRC_i_Message[138] ^ CRC_i_Message[137] ^ CRC_i_Message[133] ^ CRC_i_Message[131] ^ CRC_i_Message[130] ^ CRC_i_Message[129] ^ CRC_i_Message[128] ^ CRC_i_Message[124] ^ CRC_i_Message[122] ^ CRC_i_Message[121] ^ CRC_i_Message[120] ^ CRC_i_Message[119] ^ CRC_i_Message[113] ^ CRC_i_Message[112] ^ CRC_i_Message[107] ^ CRC_i_Message[105] ^ CRC_i_Message[101] ^ CRC_i_Message[100] ^ CRC_i_Message[98] ^ CRC_i_Message[95] ^ CRC_i_Message[94] ^ CRC_i_Message[90] ^ CRC_i_Message[89] ^ CRC_i_Message[87] ^ CRC_i_Message[86] ^ CRC_i_Message[85] ^ CRC_i_Message[84] ^ CRC_i_Message[74] ^ CRC_i_Message[73] ^ CRC_i_Message[70] ^ CRC_i_Message[68] ^ CRC_i_Message[66] ^ CRC_i_Message[65] ^ CRC_i_Message[64] ^ CRC_i_Message[63] ^ CRC_i_Message[62] ^ CRC_i_Message[59] ^ CRC_i_Message[58] ^ CRC_i_Message[57] ^ CRC_i_Message[55] ^ CRC_i_Message[54] ^ CRC_i_Message[53] ^ CRC_i_Message[49] ^ CRC_i_Message[48] ^ CRC_i_Message[47] ^ CRC_i_Message[46] ^ CRC_i_Message[44] ^ CRC_i_Message[42] ^ CRC_i_Message[40] ^ CRC_i_Message[32] ^ CRC_i_Message[30] ^ CRC_i_Message[29] ^ CRC_i_Message[28] ^ CRC_i_Message[26] ^ CRC_i_Message[22] ^ CRC_i_Message[19] ^ CRC_i_Message[13] ^ CRC_i_Message[8] ^ CRC_i_Message[4] ^ CRC_i_Message[1]);
		end	
        else begin
            CRC_o_CRC   = {POLY_WIDTH{1'b0}};
        end
    end
    else begin
        CRC_o_CRC   = {POLY_WIDTH{1'b0}};
    end
end
/* Instantiations */

endmodule
/*********** END_OF_FILE ***********/